-------------------------------------------------------------------------------
-- Title      : mux_4_1
-- Project    : 
-------------------------------------------------------------------------------
-- File       : mux_4_1.vhdl
-- Author     : Collin Clark  <collinclark@wifi-roaming-128-4-155-167.host.udel.edu>
-- Company    : 
-- Created    : 2018-03-11
-- Last update: 2018-03-11
-- Platform   : 
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description: 
-------------------------------------------------------------------------------
-- Copyright (c) 2018 
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2018-03-11  1.0      collinclark	Created
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

-------------------------------------------------------------------------------

entity mux_4_1 is

  generic (word0 : integer := 0;
           word1 : integer := 1;
           word2 : integer := 2;
           word3 : integer := 3;
           
    );

  port (switch : std_logic_vector(1 downto 0)
    );

end entity mux_4_1;

-------------------------------------------------------------------------------

architecture str of mux_4_1 is

  -----------------------------------------------------------------------------
  -- Internal signal declarations
  -----------------------------------------------------------------------------

begin  -- architecture str

  -----------------------------------------------------------------------------
  -- Component instantiations
  -----------------------------------------------------------------------------

end architecture str;

-------------------------------------------------------------------------------
